library verilog;
use verilog.vl_types.all;
entity eth_tb is
end eth_tb;
