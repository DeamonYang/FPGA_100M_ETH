library verilog;
use verilog.vl_types.all;
entity ip_proto_test_tb is
end ip_proto_test_tb;
