library verilog;
use verilog.vl_types.all;
entity udp_proto_test_tb is
end udp_proto_test_tb;
