library verilog;
use verilog.vl_types.all;
entity check_sum_tb is
end check_sum_tb;
